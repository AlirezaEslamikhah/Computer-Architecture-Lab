-- implementing a module that distinguishes 110 with type and case-when 
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
